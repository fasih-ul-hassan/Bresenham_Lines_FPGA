module Test();
	
	reg reset, clk;
	wire [7:0] x;
	wire [6:0] y;
	
	xy_coordinates UU (clk, reset, x, y);
	initial
	begin
	reset = 1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	reset = 0; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	reset = 1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	clk=0; #10; clk=1; #10;		clk=0; #10; clk=1; #10;
	end
endmodule
